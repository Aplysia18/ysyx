module ysyx_24110015_AXIArbiter (
    input clk,
    input rst

);


endmodule