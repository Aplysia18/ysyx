module ysyx_24110015_IFU (
  input clk,
  input rst,
  input [31:0] pc,
  output [31:0] inst
);


endmodule